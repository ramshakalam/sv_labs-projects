class id_entry;
    bit [3:0] id;
    bit [3:0] master_id;
    bit [3:0] slave_id;
    bit       is_read;
endclass